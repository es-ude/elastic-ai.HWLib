-- A LUT version of sigmoid
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;               -- for type conversions

entity sigmoid is
    port (
        x : in signed(15 downto 0);
        y : out signed(15 downto 0)
    );

end sigmoid;

architecture rtl of sigmoid is
begin
    
    sigmoid_process:process(x)
    begin
        if x<="1111101101000110" then
            y <= "0000000000000000"; -- 0
        elsif x<="1111110001100100" then
            y <= "0000000000000101"; -- 5
        elsif x<="1111110011100011" then
            y <= "0000000000001001"; -- 9
        elsif x<="1111110100111000" then
            y <= "0000000000001101"; -- 13
        elsif x<="1111110101111010" then
            y <= "0000000000010001"; -- 17
        elsif x<="1111110110110000" then
            y <= "0000000000010101"; -- 21
        elsif x<="1111110111011110" then
            y <= "0000000000011001"; -- 25
        elsif x<="1111111000000110" then
            y <= "0000000000011101"; -- 29
        elsif x<="1111111000101001" then
            y <= "0000000000100001"; -- 33
        elsif x<="1111111001001010" then
            y <= "0000000000100101"; -- 37
        elsif x<="1111111001101000" then
            y <= "0000000000101001"; -- 41
        elsif x<="1111111010000011" then
            y <= "0000000000101101"; -- 45
        elsif x<="1111111010011101" then
            y <= "0000000000110001"; -- 49
        elsif x<="1111111010110110" then
            y <= "0000000000110101"; -- 53
        elsif x<="1111111011001101" then
            y <= "0000000000111001"; -- 57
        elsif x<="1111111011100011" then
            y <= "0000000000111101"; -- 61
        elsif x<="1111111011111000" then
            y <= "0000000001000001"; -- 65
        elsif x<="1111111100001101" then
            y <= "0000000001000101"; -- 69
        elsif x<="1111111100100000" then
            y <= "0000000001001001"; -- 73
        elsif x<="1111111100110011" then
            y <= "0000000001001101"; -- 77
        elsif x<="1111111101000110" then
            y <= "0000000001010001"; -- 81
        elsif x<="1111111101011000" then
            y <= "0000000001010101"; -- 85
        elsif x<="1111111101101010" then
            y <= "0000000001011001"; -- 89
        elsif x<="1111111101111011" then
            y <= "0000000001011101"; -- 93
        elsif x<="1111111110001100" then
            y <= "0000000001100001"; -- 97
        elsif x<="1111111110011101" then
            y <= "0000000001100101"; -- 101
        elsif x<="1111111110101101" then
            y <= "0000000001101001"; -- 105
        elsif x<="1111111110111110" then
            y <= "0000000001101101"; -- 109
        elsif x<="1111111111001110" then
            y <= "0000000001110001"; -- 113
        elsif x<="1111111111011110" then
            y <= "0000000001110101"; -- 117
        elsif x<="1111111111101110" then
            y <= "0000000001111001"; -- 121
        elsif x<="1111111111111110" then
            y <= "0000000001111101"; -- 125
        elsif x<="0000000000001110" then
            y <= "0000000010000001"; -- 129
        elsif x<="0000000000011110" then
            y <= "0000000010000101"; -- 133
        elsif x<="0000000000101110" then
            y <= "0000000010001001"; -- 137
        elsif x<="0000000000111110" then
            y <= "0000000010001101"; -- 141
        elsif x<="0000000001001110" then
            y <= "0000000010010001"; -- 145
        elsif x<="0000000001011111" then
            y <= "0000000010010101"; -- 149
        elsif x<="0000000001110000" then
            y <= "0000000010011001"; -- 153
        elsif x<="0000000010000001" then
            y <= "0000000010011101"; -- 157
        elsif x<="0000000010010010" then
            y <= "0000000010100001"; -- 161
        elsif x<="0000000010100100" then
            y <= "0000000010100101"; -- 165
        elsif x<="0000000010110110" then
            y <= "0000000010101001"; -- 169
        elsif x<="0000000011001000" then
            y <= "0000000010101101"; -- 173
        elsif x<="0000000011011011" then
            y <= "0000000010110001"; -- 177
        elsif x<="0000000011101110" then
            y <= "0000000010110101"; -- 181
        elsif x<="0000000100000011" then
            y <= "0000000010111001"; -- 185
        elsif x<="0000000100011000" then
            y <= "0000000010111101"; -- 189
        elsif x<="0000000100101101" then
            y <= "0000000011000001"; -- 193
        elsif x<="0000000101000100" then
            y <= "0000000011000101"; -- 197
        elsif x<="0000000101011100" then
            y <= "0000000011001001"; -- 201
        elsif x<="0000000101110110" then
            y <= "0000000011001101"; -- 205
        elsif x<="0000000110010001" then
            y <= "0000000011010001"; -- 209
        elsif x<="0000000110101110" then
            y <= "0000000011010101"; -- 213
        elsif x<="0000000111001110" then
            y <= "0000000011011001"; -- 217
        elsif x<="0000000111110001" then
            y <= "0000000011011101"; -- 221
        elsif x<="0000001000011000" then
            y <= "0000000011100001"; -- 225
        elsif x<="0000001001000100" then
            y <= "0000000011100101"; -- 229
        elsif x<="0000001001111000" then
            y <= "0000000011101001"; -- 233
        elsif x<="0000001010110110" then
            y <= "0000000011101101"; -- 237
        elsif x<="0000001100000101" then
            y <= "0000000011110001"; -- 241
        elsif x<="0000001101110110" then
            y <= "0000000011110101"; -- 245
        elsif x<="0000010001001001" then
            y <= "0000000011111001"; -- 249
        else
            y <= "0000000100000000"; -- 256
        end if;
    end process;
end rtl;


