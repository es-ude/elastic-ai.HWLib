-- A LUT version of tanh
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;               -- for type conversions

entity tanh is
    port (
        x : in signed(15 downto 0);
        y : out signed(15 downto 0)
    );

end tanh;

architecture rtl of tanh is
begin
    
    tanh_process:process(x)
    begin
        if x<="1111110110100100" then
            y <= "1111111100000000"; -- -256
        elsif x<="1111111000110011" then
            y <= "1111111100010011"; -- -237
        elsif x<="1111111001110010" then
            y <= "1111111100011011"; -- -229
        elsif x<="1111111010011101" then
            y <= "1111111100100011"; -- -221
        elsif x<="1111111010111110" then
            y <= "1111111100101011"; -- -213
        elsif x<="1111111011011001" then
            y <= "1111111100110011"; -- -205
        elsif x<="1111111011110000" then
            y <= "1111111100111011"; -- -197
        elsif x<="1111111100000100" then
            y <= "1111111101000011"; -- -189
        elsif x<="1111111100010110" then
            y <= "1111111101001011"; -- -181
        elsif x<="1111111100100110" then
            y <= "1111111101010011"; -- -173
        elsif x<="1111111100110101" then
            y <= "1111111101011011"; -- -165
        elsif x<="1111111101000011" then
            y <= "1111111101100011"; -- -157
        elsif x<="1111111101010000" then
            y <= "1111111101101100"; -- -148
        elsif x<="1111111101011100" then
            y <= "1111111101110100"; -- -140
        elsif x<="1111111101101000" then
            y <= "1111111101111100"; -- -132
        elsif x<="1111111101110011" then
            y <= "1111111110000100"; -- -124
        elsif x<="1111111101111101" then
            y <= "1111111110001100"; -- -116
        elsif x<="1111111110001000" then
            y <= "1111111110010100"; -- -108
        elsif x<="1111111110010001" then
            y <= "1111111110011100"; -- -100
        elsif x<="1111111110011011" then
            y <= "1111111110100100"; -- -92
        elsif x<="1111111110100100" then
            y <= "1111111110101100"; -- -84
        elsif x<="1111111110101101" then
            y <= "1111111110110100"; -- -76
        elsif x<="1111111110110110" then
            y <= "1111111110111100"; -- -68
        elsif x<="1111111110111111" then
            y <= "1111111111000100"; -- -60
        elsif x<="1111111111001000" then
            y <= "1111111111001100"; -- -52
        elsif x<="1111111111010000" then
            y <= "1111111111010101"; -- -43
        elsif x<="1111111111011000" then
            y <= "1111111111011101"; -- -35
        elsif x<="1111111111100001" then
            y <= "1111111111100101"; -- -27
        elsif x<="1111111111101001" then
            y <= "1111111111101101"; -- -19
        elsif x<="1111111111110001" then
            y <= "1111111111110101"; -- -11
        elsif x<="1111111111111001" then
            y <= "1111111111111101"; -- -3
        elsif x<="0000000000000000" then
            y <= "0000000000000100"; -- 4
        elsif x<="0000000000001000" then
            y <= "0000000000001100"; -- 12
        elsif x<="0000000000010000" then
            y <= "0000000000010100"; -- 20
        elsif x<="0000000000011000" then
            y <= "0000000000011100"; -- 28
        elsif x<="0000000000100001" then
            y <= "0000000000100100"; -- 36
        elsif x<="0000000000101001" then
            y <= "0000000000101100"; -- 44
        elsif x<="0000000000110001" then
            y <= "0000000000110101"; -- 53
        elsif x<="0000000000111010" then
            y <= "0000000000111101"; -- 61
        elsif x<="0000000001000010" then
            y <= "0000000001000101"; -- 69
        elsif x<="0000000001001011" then
            y <= "0000000001001101"; -- 77
        elsif x<="0000000001010100" then
            y <= "0000000001010101"; -- 85
        elsif x<="0000000001011101" then
            y <= "0000000001011101"; -- 93
        elsif x<="0000000001100110" then
            y <= "0000000001100101"; -- 101
        elsif x<="0000000001110000" then
            y <= "0000000001101101"; -- 109
        elsif x<="0000000001111010" then
            y <= "0000000001110101"; -- 117
        elsif x<="0000000010000100" then
            y <= "0000000001111101"; -- 125
        elsif x<="0000000010001111" then
            y <= "0000000010000101"; -- 133
        elsif x<="0000000010011010" then
            y <= "0000000010001101"; -- 141
        elsif x<="0000000010100101" then
            y <= "0000000010010101"; -- 149
        elsif x<="0000000010110010" then
            y <= "0000000010011110"; -- 158
        elsif x<="0000000010111111" then
            y <= "0000000010100110"; -- 166
        elsif x<="0000000011001101" then
            y <= "0000000010101110"; -- 174
        elsif x<="0000000011011100" then
            y <= "0000000010110110"; -- 182
        elsif x<="0000000011101100" then
            y <= "0000000010111110"; -- 190
        elsif x<="0000000011111110" then
            y <= "0000000011000110"; -- 198
        elsif x<="0000000100010011" then
            y <= "0000000011001110"; -- 206
        elsif x<="0000000100101010" then
            y <= "0000000011010110"; -- 214
        elsif x<="0000000101000110" then
            y <= "0000000011011110"; -- 222
        elsif x<="0000000101100111" then
            y <= "0000000011100110"; -- 230
        elsif x<="0000000110010100" then
            y <= "0000000011101110"; -- 238
        elsif x<="0000000111011000" then
            y <= "0000000011110110"; -- 246
        elsif x<="0000001010010000" then
            y <= "0000000011111111"; -- 255
        else
            y <= "0000000100000000"; -- 256
        end if;
    end process;
end rtl;